clkpll_inst : clkpll PORT MAP (
		inclk0	 => inclk0_sig,
		c0	 => c0_sig,
		locked	 => locked_sig
	);
